// 讓output 永遠等於1

module top_module( output one );
	
	assign one = 1'b1;
endmodule